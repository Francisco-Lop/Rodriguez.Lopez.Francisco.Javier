** Profile: "SCHEMATIC1-rectificacion-en-puente-practica3"  [ C:\Users\emile\Desktop\practica 3 garabito\rectificador monofasico en puente practica 3-pspicefiles\schematic1\rectificacion-en-puente-practica3.sim ] 

** Creating circuit file "rectificacion-en-puente-practica3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60ms 0 10ms 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
