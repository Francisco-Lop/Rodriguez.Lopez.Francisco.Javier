** Profile: "SCHEMATIC1-fourier"  [ C:\Cadence\SPB_16.5\tools\capture\parte 2,1-pspicefiles\schematic1\fourier.sim ] 

** Creating circuit file "fourier.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN 10us 60ms 10ms 60ms SKIPBP 
.FOUR 60 2 1 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
